module Spartan6_DSP48A1(A,B,D,C,CLK,CARRYIN,OPMODE,BCIN,RSTA,RSTB,RSTM,RSTP,RSTC,RSTD,RSTCARRYIN,RSTOPMODE,CEA,CEB,CEM,CEP,CEC,CED,CECARRYIN,CEOPMODE,PCIN,BCOUT,PCOUT,P,M,CARRYOUT,CARRYOUTF);
//Parameters
parameter A0REG=1'b0;
parameter A1REG=1'b1;
parameter B0REG=1'b0;
parameter B1REG=1'b1;
parameter CREG=1'b1;
parameter DREG=1'b1;
parameter MREG=1'b1;
parameter PREG=1'b1;
parameter CARRTINREG=1'b1;
parameter CARRYOUTREG=1'b1;
parameter OPMODEREG=1'b1;
parameter CARRYINSEL="OPMODE5";//or CARRYIN if it is input of user or if it is none the output of mux is 0
parameter B_INPUT="DIRECT";//or CASCADE if it is from BCIN as input or if it is none the output of mux is 0
parameter RSTTYPE="SYNC";//or ASYNE if it is asynchronus

//Data Ports
input [17:0]A;
input [17:0]B;
input [17:0]BCIN;
input [47:0]C;
input [17:0]D;
input CARRYIN;
output [35:0]M;
output [47:0]P;
output CARRYOUT;
output CARRYOUTF;
//Control Input Ports
input CLK;
input [7:0]OPMODE;
//Clock Enable Input Ports
input CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP;
//Reset Input Ports
input RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP;
//Cascade Ports
input [47:0]PCIN;
output [17:0]BCOUT;
output[47:0]PCOUT;
//Wires
wire [17:0] D_WIRE;
wire [17:0] B_IN_WIRE;
wire [17:0] B0_WIRE;
wire [17:0] B1_WIRE;
wire [17:0] A0_WIRE;
wire [17:0] A1_WIRE;
wire [47:0] C_WIRE;
wire [35:0] M_WIRE;
wire [47:0] P_WIRE;
wire [17:0] D_B0_WIRE;
wire [17:0] D_B0_MUX_WIRE;
wire [35:0] A1_B1_WIRE;
wire [47:0] D_A_B_WIRE;
wire [47:0] X_MUX_WIRE;
wire [47:0] Z_MUX_WIRE;
wire [47:0] X_Z_WIRE;
wire [7:0] OPMODE_WIRE;
wire CARRYIN_WIRE;
wire CYI_WIRE;
wire CARRYOUT_WIRE;
wire CYO_WIRE;
//Instantiations
REG_MUX #(18,RSTTYPE) REG_D(.INPUT(D),.SEL(DREG[0]),.RST(RSTD),.CLK(CLK),.CE(CED),.OUTPUT(D_WIRE));
REG_MUX #(18,RSTTYPE) RGE_B0(.INPUT(B_IN_WIRE),.SEL(B0REG[0]),.RST(RSTB),.CLK(CLK),.CE(CEB),.OUTPUT(B0_WIRE));
REG_MUX #(18,RSTTYPE) REG_A0(.INPUT(A),.SEL(A0REG[0]),.RST(RSTA),.CLK(CLK),.CE(CEA),.OUTPUT(A0_WIRE));
REG_MUX #(48,RSTTYPE) REG_C(.INPUT(C),.SEL(CREG[0]),.RST(RSTC),.CLK(CLK),.CE(CEC),.OUTPUT(C_WIRE));
REG_MUX #(18,RSTTYPE) RGE_B1(.INPUT(D_B0_MUX_WIRE),.SEL(B1REG[0]),.RST(RSTB),.CLK(CLK),.CE(CEB),.OUTPUT(B1_WIRE));
REG_MUX #(18,RSTTYPE) REG_A1(.INPUT(A0_WIRE),.SEL(A1REG[0]),.RST(RSTA),.CLK(CLK),.CE(CEA),.OUTPUT(A1_WIRE));
REG_MUX #(36,RSTTYPE) REG_M(.INPUT(A1_B1_WIRE),.SEL(MREG[0]),.RST(RSTM),.CLK(CLK),.CE(CEM),.OUTPUT(M_WIRE));
REG_MUX #(48,RSTTYPE) REG_P(.INPUT(X_Z_WIRE),.SEL(PREG[0]),.RST(RSTP),.CLK(CLK),.CE(CEP),.OUTPUT(P_WIRE));
REG_MUX #(8,RSTTYPE) REG_OPMODE(.INPUT(OPMODE),.SEL(OPMODEREG[0]),.RST(RSTOPMODE),.CLK(CLK),.CE(CEOPMODE),.OUTPUT(OPMODE_WIRE));
REG_MUX #(1,RSTTYPE) CYI(.INPUT(CARRYIN_WIRE),.SEL(CARRTINREG[0]),.RST(RSTCARRYIN),.CLK(CLK),.CE(CECARRYIN),.OUTPUT(CYI_WIRE));
REG_MUX #(1,RSTTYPE) CYO(.INPUT(CARRYOUT_WIRE),.SEL(CARRYOUTREG[0]),.RST(1'b0),.CLK(CLK),.CE(1'b0),.OUTPUT(CYO_WIRE));


MUX_4_1 #(48) MUX_X(.IN0(D_A_B_WIRE),.IN1(P_WIRE),.IN2({12'h000,M_WIRE}),.IN3(48'h000000000000),.SEL(OPMODE_WIRE[1:0]),.OUT(X_MUX_WIRE));
MUX_4_1 #(48) MUX_Z(.IN0(C_WIRE),.IN1(P_WIRE),.IN2(PCIN),.IN3(48'h000000000000),.SEL(OPMODE_WIRE[3:2]),.OUT(Z_MUX_WIRE));

assign B_IN_WIRE=(B_INPUT=="DIRECT")?B:(B_INPUT=="CASCADE")?BCIN:0;
assign D_B0_WIRE=(OPMODE_WIRE[6])?(D_WIRE-B0_WIRE):(D_WIRE+B0_WIRE);
assign D_B0_MUX_WIRE=(OPMODE_WIRE[4])?D_B0_WIRE:B0_WIRE;
assign A1_B1_WIRE=A1_WIRE*B1_WIRE;
assign D_A_B_WIRE={D_WIRE[11:0],A1_WIRE,B1_WIRE};
assign M=M_WIRE;
assign BCOUT=B1_WIRE;
assign CARRYIN_WIRE=(CARRYINSEL=="OPMODE5")?OPMODE_WIRE[5]:(CARRYINSEL=="CARRYIN")?CARRYIN:0;
assign{CARRYOUT_WIRE,X_Z_WIRE}=(OPMODE_WIRE[7])?Z_MUX_WIRE-(X_MUX_WIRE+CYI_WIRE) :X_MUX_WIRE+Z_MUX_WIRE+CYI_WIRE;
assign P=P_WIRE;
assign PCOUT=P_WIRE;
assign CARRYOUT=CYO_WIRE;
assign CARRYOUTF=CYO_WIRE;

endmodule
